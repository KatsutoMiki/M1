`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/01/27 13:55:18
// Design Name: 
// Module Name: dfil_new_reg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dfil_new_reg(
        input wire indata,
        input CLK,
        output wire [29:0] sum,
        output wire out
    );

    reg [14:0] count_pulse = 15'b0;
    reg [14:0] clk_counter = 15'd0;
    reg [4999:0] filter=0;
    reg fil= 1'b0;
    reg [29:0] reg_sum = 30'b0;
    // reg [15:0] new_result = 0;
    // reg [15:0] old_result = 0;
    reg state = 0;
    reg full = 0;
    parameter STACK = 0;
    parameter WATING = 1;
    parameter GENERATE_PULSE = 2;
    parameter WATING_TIME = 16'd0;
    parameter WATING_SUM = 5'b11111;

    always@(posedge CLK)begin

        filter <= {filter[4999:0], indata};

         // if (state) begin
        //     if (filter[0] == 1 & filter[4999] == 0) begin
        //         reg_sum <= reg_sum + 1;    
        //     end
        //     else if (filter[0] == 0 & filter[4999] == 1) begin
        //         reg_sum <= reg_sum - 1;
        //     end
        //     else begin
        //         reg_sum <= reg_sum;
        //     end

        //     if(reg_sum > 14'd4500)begin
        //         fil <= 1'b1;
        //     end
        //     if(reg_sum < 14'd500)begin
        //         fil <= 1'b0;
        //     end
        // end
        // else begin
        //     clk_counter <= clk_counter + 1;
        //     if (clk_counter == WATING_TIME)begin
        //         state <= 1;
        //     end
        // end
		count_pulse <= filter[0]+filter[1]+filter[2]+filter[3]+filter[4]+filter[5]+filter[6]+filter[7]+filter[8]+filter[9]+filter[10]+filter[11]+filter[12]+filter[13]+filter[14]+filter[15]+filter[16]+filter[17]+filter[18]+filter[19]+filter[20]+filter[21]+filter[22]+filter[23]+filter[24]+filter[25]+filter[26]+filter[27]+filter[28]+filter[29]+filter[30]+filter[31]+filter[32]+filter[33]+filter[34]+filter[35]+filter[36]+filter[37]+filter[38]+filter[39]+filter[40]+filter[41]+filter[42]+filter[43]+filter[44]+filter[45]+filter[46]+filter[47]+filter[48]+filter[49]+filter[50]+filter[51]+filter[52]+filter[53]+filter[54]+filter[55]+filter[56]+filter[57]+filter[58]+filter[59]+filter[60]+filter[61]+filter[62]+filter[63]+filter[64]+filter[65]+filter[66]+filter[67]+filter[68]+filter[69]+filter[70]+filter[71]+filter[72]+filter[73]+filter[74]+filter[75]+filter[76]+filter[77]+filter[78]+filter[79]+filter[80]+filter[81]+filter[82]+filter[83]+filter[84]+filter[85]+filter[86]+filter[87]+filter[88]+filter[89]+filter[90]+filter[91]+filter[92]+filter[93]+filter[94]+filter[95]+filter[96]+filter[97]+filter[98]+filter[99]+filter[100]+filter[101]+filter[102]+filter[103]+filter[104]+filter[105]+filter[106]+filter[107]+filter[108]+filter[109]+filter[110]+filter[111]+filter[112]+filter[113]+filter[114]+filter[115]+filter[116]+filter[117]+filter[118]+filter[119]+filter[120]+filter[121]+filter[122]+filter[123]+filter[124]+filter[125]+filter[126]+filter[127]+filter[128]+filter[129]+filter[130]+filter[131]+filter[132]+filter[133]+filter[134]+filter[135]+filter[136]+filter[137]+filter[138]+filter[139]+filter[140]+filter[141]+filter[142]+filter[143]+filter[144]+filter[145]+filter[146]+filter[147]+filter[148]+filter[149]+filter[150]+filter[151]+filter[152]+filter[153]+filter[154]+filter[155]+filter[156]+filter[157]+filter[158]+filter[159]+filter[160]+filter[161]+filter[162]+filter[163]+filter[164]+filter[165]+filter[166]+filter[167]+filter[168]+filter[169]+filter[170]+filter[171]+filter[172]+filter[173]+filter[174]+filter[175]+filter[176]+filter[177]+filter[178]+filter[179]+filter[180]+filter[181]+filter[182]+filter[183]+filter[184]+filter[185]+filter[186]+filter[187]+filter[188]+filter[189]+filter[190]+filter[191]+filter[192]+filter[193]+filter[194]+filter[195]+filter[196]+filter[197]+filter[198]+filter[199]+filter[200]+filter[201]+filter[202]+filter[203]+filter[204]+filter[205]+filter[206]+filter[207]+filter[208]+filter[209]+filter[210]+filter[211]+filter[212]+filter[213]+filter[214]+filter[215]+filter[216]+filter[217]+filter[218]+filter[219]+filter[220]+filter[221]+filter[222]+filter[223]+filter[224]+filter[225]+filter[226]+filter[227]+filter[228]+filter[229]+filter[230]+filter[231]+filter[232]+filter[233]+filter[234]+filter[235]+filter[236]+filter[237]+filter[238]+filter[239]+filter[240]+filter[241]+filter[242]+filter[243]+filter[244]+filter[245]+filter[246]+filter[247]+filter[248]+filter[249]+filter[250]+filter[251]+filter[252]+filter[253]+filter[254]+filter[255]+filter[256]+filter[257]+filter[258]+filter[259]+filter[260]+filter[261]+filter[262]+filter[263]+filter[264]+filter[265]+filter[266]+filter[267]+filter[268]+filter[269]+filter[270]+filter[271]+filter[272]+filter[273]+filter[274]+filter[275]+filter[276]+filter[277]+filter[278]+filter[279]+filter[280]+filter[281]+filter[282]+filter[283]+filter[284]+filter[285]+filter[286]+filter[287]+filter[288]+filter[289]+filter[290]+filter[291]+filter[292]+filter[293]+filter[294]+filter[295]+filter[296]+filter[297]+filter[298]+filter[299]+filter[300]+filter[301]+filter[302]+filter[303]+filter[304]+filter[305]+filter[306]+filter[307]+filter[308]+filter[309]+filter[310]+filter[311]+filter[312]+filter[313]+filter[314]+filter[315]+filter[316]+filter[317]+filter[318]+filter[319]+filter[320]+filter[321]+filter[322]+filter[323]+filter[324]+filter[325]+filter[326]+filter[327]+filter[328]+filter[329]+filter[330]+filter[331]+filter[332]+filter[333]+filter[334]+filter[335]+filter[336]+filter[337]+filter[338]+filter[339]+filter[340]+filter[341]+filter[342]+filter[343]+filter[344]+filter[345]+filter[346]+filter[347]+filter[348]+filter[349]+filter[350]+filter[351]+filter[352]+filter[353]+filter[354]+filter[355]+filter[356]+filter[357]+filter[358]+filter[359]+filter[360]+filter[361]+filter[362]+filter[363]+filter[364]+filter[365]+filter[366]+filter[367]+filter[368]+filter[369]+filter[370]+filter[371]+filter[372]+filter[373]+filter[374]+filter[375]+filter[376]+filter[377]+filter[378]+filter[379]+filter[380]+filter[381]+filter[382]+filter[383]+filter[384]+filter[385]+filter[386]+filter[387]+filter[388]+filter[389]+filter[390]+filter[391]+filter[392]+filter[393]+filter[394]+filter[395]+filter[396]+filter[397]+filter[398]+filter[399]+filter[400]+filter[401]+filter[402]+filter[403]+filter[404]+filter[405]+filter[406]+filter[407]+filter[408]+filter[409]+filter[410]+filter[411]+filter[412]+filter[413]+filter[414]+filter[415]+filter[416]+filter[417]+filter[418]+filter[419]+filter[420]+filter[421]+filter[422]+filter[423]+filter[424]+filter[425]+filter[426]+filter[427]+filter[428]+filter[429]+filter[430]+filter[431]+filter[432]+filter[433]+filter[434]+filter[435]+filter[436]+filter[437]+filter[438]+filter[439]+filter[440]+filter[441]+filter[442]+filter[443]+filter[444]+filter[445]+filter[446]+filter[447]+filter[448]+filter[449]+filter[450]+filter[451]+filter[452]+filter[453]+filter[454]+filter[455]+filter[456]+filter[457]+filter[458]+filter[459]+filter[460]+filter[461]+filter[462]+filter[463]+filter[464]+filter[465]+filter[466]+filter[467]+filter[468]+filter[469]+filter[470]+filter[471]+filter[472]+filter[473]+filter[474]+filter[475]+filter[476]+filter[477]+filter[478]+filter[479]+filter[480]+filter[481]+filter[482]+filter[483]+filter[484]+filter[485]+filter[486]+filter[487]+filter[488]+filter[489]+filter[490]+filter[491]+filter[492]+filter[493]+filter[494]+filter[495]+filter[496]+filter[497]+filter[498]+filter[499]+filter[500]+filter[501]+filter[502]+filter[503]+filter[504]+filter[505]+filter[506]+filter[507]+filter[508]+filter[509]+filter[510]+filter[511]+filter[512]+filter[513]+filter[514]+filter[515]+filter[516]+filter[517]+filter[518]+filter[519]+filter[520]+filter[521]+filter[522]+filter[523]+filter[524]+filter[525]+filter[526]+filter[527]+filter[528]+filter[529]+filter[530]+filter[531]+filter[532]+filter[533]+filter[534]+filter[535]+filter[536]+filter[537]+filter[538]+filter[539]+filter[540]+filter[541]+filter[542]+filter[543]+filter[544]+filter[545]+filter[546]+filter[547]+filter[548]+filter[549]+filter[550]+filter[551]+filter[552]+filter[553]+filter[554]+filter[555]+filter[556]+filter[557]+filter[558]+filter[559]+filter[560]+filter[561]+filter[562]+filter[563]+filter[564]+filter[565]+filter[566]+filter[567]+filter[568]+filter[569]+filter[570]+filter[571]+filter[572]+filter[573]+filter[574]+filter[575]+filter[576]+filter[577]+filter[578]+filter[579]+filter[580]+filter[581]+filter[582]+filter[583]+filter[584]+filter[585]+filter[586]+filter[587]+filter[588]+filter[589]+filter[590]+filter[591]+filter[592]+filter[593]+filter[594]+filter[595]+filter[596]+filter[597]+filter[598]+filter[599]+filter[600]+filter[601]+filter[602]+filter[603]+filter[604]+filter[605]+filter[606]+filter[607]+filter[608]+filter[609]+filter[610]+filter[611]+filter[612]+filter[613]+filter[614]+filter[615]+filter[616]+filter[617]+filter[618]+filter[619]+filter[620]+filter[621]+filter[622]+filter[623]+filter[624]+filter[625]+filter[626]+filter[627]+filter[628]+filter[629]+filter[630]+filter[631]+filter[632]+filter[633]+filter[634]+filter[635]+filter[636]+filter[637]+filter[638]+filter[639]+filter[640]+filter[641]+filter[642]+filter[643]+filter[644]+filter[645]+filter[646]+filter[647]+filter[648]+filter[649]+filter[650]+filter[651]+filter[652]+filter[653]+filter[654]+filter[655]+filter[656]+filter[657]+filter[658]+filter[659]+filter[660]+filter[661]+filter[662]+filter[663]+filter[664]+filter[665]+filter[666]+filter[667]+filter[668]+filter[669]+filter[670]+filter[671]+filter[672]+filter[673]+filter[674]+filter[675]+filter[676]+filter[677]+filter[678]+filter[679]+filter[680]+filter[681]+filter[682]+filter[683]+filter[684]+filter[685]+filter[686]+filter[687]+filter[688]+filter[689]+filter[690]+filter[691]+filter[692]+filter[693]+filter[694]+filter[695]+filter[696]+filter[697]+filter[698]+filter[699]+filter[700]+filter[701]+filter[702]+filter[703]+filter[704]+filter[705]+filter[706]+filter[707]+filter[708]+filter[709]+filter[710]+filter[711]+filter[712]+filter[713]+filter[714]+filter[715]+filter[716]+filter[717]+filter[718]+filter[719]+filter[720]+filter[721]+filter[722]+filter[723]+filter[724]+filter[725]+filter[726]+filter[727]+filter[728]+filter[729]+filter[730]+filter[731]+filter[732]+filter[733]+filter[734]+filter[735]+filter[736]+filter[737]+filter[738]+filter[739]+filter[740]+filter[741]+filter[742]+filter[743]+filter[744]+filter[745]+filter[746]+filter[747]+filter[748]+filter[749]+filter[750]+filter[751]+filter[752]+filter[753]+filter[754]+filter[755]+filter[756]+filter[757]+filter[758]+filter[759]+filter[760]+filter[761]+filter[762]+filter[763]+filter[764]+filter[765]+filter[766]+filter[767]+filter[768]+filter[769]+filter[770]+filter[771]+filter[772]+filter[773]+filter[774]+filter[775]+filter[776]+filter[777]+filter[778]+filter[779]+filter[780]+filter[781]+filter[782]+filter[783]+filter[784]+filter[785]+filter[786]+filter[787]+filter[788]+filter[789]+filter[790]+filter[791]+filter[792]+filter[793]+filter[794]+filter[795]+filter[796]+filter[797]+filter[798]+filter[799]+filter[800]+filter[801]+filter[802]+filter[803]+filter[804]+filter[805]+filter[806]+filter[807]+filter[808]+filter[809]+filter[810]+filter[811]+filter[812]+filter[813]+filter[814]+filter[815]+filter[816]+filter[817]+filter[818]+filter[819]+filter[820]+filter[821]+filter[822]+filter[823]+filter[824]+filter[825]+filter[826]+filter[827]+filter[828]+filter[829]+filter[830]+filter[831]+filter[832]+filter[833]+filter[834]+filter[835]+filter[836]+filter[837]+filter[838]+filter[839]+filter[840]+filter[841]+filter[842]+filter[843]+filter[844]+filter[845]+filter[846]+filter[847]+filter[848]+filter[849]+filter[850]+filter[851]+filter[852]+filter[853]+filter[854]+filter[855]+filter[856]+filter[857]+filter[858]+filter[859]+filter[860]+filter[861]+filter[862]+filter[863]+filter[864]+filter[865]+filter[866]+filter[867]+filter[868]+filter[869]+filter[870]+filter[871]+filter[872]+filter[873]+filter[874]+filter[875]+filter[876]+filter[877]+filter[878]+filter[879]+filter[880]+filter[881]+filter[882]+filter[883]+filter[884]+filter[885]+filter[886]+filter[887]+filter[888]+filter[889]+filter[890]+filter[891]+filter[892]+filter[893]+filter[894]+filter[895]+filter[896]+filter[897]+filter[898]+filter[899]+filter[900]+filter[901]+filter[902]+filter[903]+filter[904]+filter[905]+filter[906]+filter[907]+filter[908]+filter[909]+filter[910]+filter[911]+filter[912]+filter[913]+filter[914]+filter[915]+filter[916]+filter[917]+filter[918]+filter[919]+filter[920]+filter[921]+filter[922]+filter[923]+filter[924]+filter[925]+filter[926]+filter[927]+filter[928]+filter[929]+filter[930]+filter[931]+filter[932]+filter[933]+filter[934]+filter[935]+filter[936]+filter[937]+filter[938]+filter[939]+filter[940]+filter[941]+filter[942]+filter[943]+filter[944]+filter[945]+filter[946]+filter[947]+filter[948]+filter[949]+filter[950]+filter[951]+filter[952]+filter[953]+filter[954]+filter[955]+filter[956]+filter[957]+filter[958]+filter[959]+filter[960]+filter[961]+filter[962]+filter[963]+filter[964]+filter[965]+filter[966]+filter[967]+filter[968]+filter[969]+filter[970]+filter[971]+filter[972]+filter[973]+filter[974]+filter[975]+filter[976]+filter[977]+filter[978]+filter[979]+filter[980]+filter[981]+filter[982]+filter[983]+filter[984]+filter[985]+filter[986]+filter[987]+filter[988]+filter[989]+filter[990]+filter[991]+filter[992]+filter[993]+filter[994]+filter[995]+filter[996]+filter[997]+filter[998]+filter[999]+filter[1000]+filter[1001]+filter[1002]+filter[1003]+filter[1004]+filter[1005]+filter[1006]+filter[1007]+filter[1008]+filter[1009]+filter[1010]+filter[1011]+filter[1012]+filter[1013]+filter[1014]+filter[1015]+filter[1016]+filter[1017]+filter[1018]+filter[1019]+filter[1020]+filter[1021]+filter[1022]+filter[1023]+filter[1024]+filter[1025]+filter[1026]+filter[1027]+filter[1028]+filter[1029]+filter[1030]+filter[1031]+filter[1032]+filter[1033]+filter[1034]+filter[1035]+filter[1036]+filter[1037]+filter[1038]+filter[1039]+filter[1040]+filter[1041]+filter[1042]+filter[1043]+filter[1044]+filter[1045]+filter[1046]+filter[1047]+filter[1048]+filter[1049]+filter[1050]+filter[1051]+filter[1052]+filter[1053]+filter[1054]+filter[1055]+filter[1056]+filter[1057]+filter[1058]+filter[1059]+filter[1060]+filter[1061]+filter[1062]+filter[1063]+filter[1064]+filter[1065]+filter[1066]+filter[1067]+filter[1068]+filter[1069]+filter[1070]+filter[1071]+filter[1072]+filter[1073]+filter[1074]+filter[1075]+filter[1076]+filter[1077]+filter[1078]+filter[1079]+filter[1080]+filter[1081]+filter[1082]+filter[1083]+filter[1084]+filter[1085]+filter[1086]+filter[1087]+filter[1088]+filter[1089]+filter[1090]+filter[1091]+filter[1092]+filter[1093]+filter[1094]+filter[1095]+filter[1096]+filter[1097]+filter[1098]+filter[1099]+filter[1100]+filter[1101]+filter[1102]+filter[1103]+filter[1104]+filter[1105]+filter[1106]+filter[1107]+filter[1108]+filter[1109]+filter[1110]+filter[1111]+filter[1112]+filter[1113]+filter[1114]+filter[1115]+filter[1116]+filter[1117]+filter[1118]+filter[1119]+filter[1120]+filter[1121]+filter[1122]+filter[1123]+filter[1124]+filter[1125]+filter[1126]+filter[1127]+filter[1128]+filter[1129]+filter[1130]+filter[1131]+filter[1132]+filter[1133]+filter[1134]+filter[1135]+filter[1136]+filter[1137]+filter[1138]+filter[1139]+filter[1140]+filter[1141]+filter[1142]+filter[1143]+filter[1144]+filter[1145]+filter[1146]+filter[1147]+filter[1148]+filter[1149]+filter[1150]+filter[1151]+filter[1152]+filter[1153]+filter[1154]+filter[1155]+filter[1156]+filter[1157]+filter[1158]+filter[1159]+filter[1160]+filter[1161]+filter[1162]+filter[1163]+filter[1164]+filter[1165]+filter[1166]+filter[1167]+filter[1168]+filter[1169]+filter[1170]+filter[1171]+filter[1172]+filter[1173]+filter[1174]+filter[1175]+filter[1176]+filter[1177]+filter[1178]+filter[1179]+filter[1180]+filter[1181]+filter[1182]+filter[1183]+filter[1184]+filter[1185]+filter[1186]+filter[1187]+filter[1188]+filter[1189]+filter[1190]+filter[1191]+filter[1192]+filter[1193]+filter[1194]+filter[1195]+filter[1196]+filter[1197]+filter[1198]+filter[1199]+filter[1200]+filter[1201]+filter[1202]+filter[1203]+filter[1204]+filter[1205]+filter[1206]+filter[1207]+filter[1208]+filter[1209]+filter[1210]+filter[1211]+filter[1212]+filter[1213]+filter[1214]+filter[1215]+filter[1216]+filter[1217]+filter[1218]+filter[1219]+filter[1220]+filter[1221]+filter[1222]+filter[1223]+filter[1224]+filter[1225]+filter[1226]+filter[1227]+filter[1228]+filter[1229]+filter[1230]+filter[1231]+filter[1232]+filter[1233]+filter[1234]+filter[1235]+filter[1236]+filter[1237]+filter[1238]+filter[1239]+filter[1240]+filter[1241]+filter[1242]+filter[1243]+filter[1244]+filter[1245]+filter[1246]+filter[1247]+filter[1248]+filter[1249]+filter[1250]+filter[1251]+filter[1252]+filter[1253]+filter[1254]+filter[1255]+filter[1256]+filter[1257]+filter[1258]+filter[1259]+filter[1260]+filter[1261]+filter[1262]+filter[1263]+filter[1264]+filter[1265]+filter[1266]+filter[1267]+filter[1268]+filter[1269]+filter[1270]+filter[1271]+filter[1272]+filter[1273]+filter[1274]+filter[1275]+filter[1276]+filter[1277]+filter[1278]+filter[1279]+filter[1280]+filter[1281]+filter[1282]+filter[1283]+filter[1284]+filter[1285]+filter[1286]+filter[1287]+filter[1288]+filter[1289]+filter[1290]+filter[1291]+filter[1292]+filter[1293]+filter[1294]+filter[1295]+filter[1296]+filter[1297]+filter[1298]+filter[1299]+filter[1300]+filter[1301]+filter[1302]+filter[1303]+filter[1304]+filter[1305]+filter[1306]+filter[1307]+filter[1308]+filter[1309]+filter[1310]+filter[1311]+filter[1312]+filter[1313]+filter[1314]+filter[1315]+filter[1316]+filter[1317]+filter[1318]+filter[1319]+filter[1320]+filter[1321]+filter[1322]+filter[1323]+filter[1324]+filter[1325]+filter[1326]+filter[1327]+filter[1328]+filter[1329]+filter[1330]+filter[1331]+filter[1332]+filter[1333]+filter[1334]+filter[1335]+filter[1336]+filter[1337]+filter[1338]+filter[1339]+filter[1340]+filter[1341]+filter[1342]+filter[1343]+filter[1344]+filter[1345]+filter[1346]+filter[1347]+filter[1348]+filter[1349]+filter[1350]+filter[1351]+filter[1352]+filter[1353]+filter[1354]+filter[1355]+filter[1356]+filter[1357]+filter[1358]+filter[1359]+filter[1360]+filter[1361]+filter[1362]+filter[1363]+filter[1364]+filter[1365]+filter[1366]+filter[1367]+filter[1368]+filter[1369]+filter[1370]+filter[1371]+filter[1372]+filter[1373]+filter[1374]+filter[1375]+filter[1376]+filter[1377]+filter[1378]+filter[1379]+filter[1380]+filter[1381]+filter[1382]+filter[1383]+filter[1384]+filter[1385]+filter[1386]+filter[1387]+filter[1388]+filter[1389]+filter[1390]+filter[1391]+filter[1392]+filter[1393]+filter[1394]+filter[1395]+filter[1396]+filter[1397]+filter[1398]+filter[1399]+filter[1400]+filter[1401]+filter[1402]+filter[1403]+filter[1404]+filter[1405]+filter[1406]+filter[1407]+filter[1408]+filter[1409]+filter[1410]+filter[1411]+filter[1412]+filter[1413]+filter[1414]+filter[1415]+filter[1416]+filter[1417]+filter[1418]+filter[1419]+filter[1420]+filter[1421]+filter[1422]+filter[1423]+filter[1424]+filter[1425]+filter[1426]+filter[1427]+filter[1428]+filter[1429]+filter[1430]+filter[1431]+filter[1432]+filter[1433]+filter[1434]+filter[1435]+filter[1436]+filter[1437]+filter[1438]+filter[1439]+filter[1440]+filter[1441]+filter[1442]+filter[1443]+filter[1444]+filter[1445]+filter[1446]+filter[1447]+filter[1448]+filter[1449]+filter[1450]+filter[1451]+filter[1452]+filter[1453]+filter[1454]+filter[1455]+filter[1456]+filter[1457]+filter[1458]+filter[1459]+filter[1460]+filter[1461]+filter[1462]+filter[1463]+filter[1464]+filter[1465]+filter[1466]+filter[1467]+filter[1468]+filter[1469]+filter[1470]+filter[1471]+filter[1472]+filter[1473]+filter[1474]+filter[1475]+filter[1476]+filter[1477]+filter[1478]+filter[1479]+filter[1480]+filter[1481]+filter[1482]+filter[1483]+filter[1484]+filter[1485]+filter[1486]+filter[1487]+filter[1488]+filter[1489]+filter[1490]+filter[1491]+filter[1492]+filter[1493]+filter[1494]+filter[1495]+filter[1496]+filter[1497]+filter[1498]+filter[1499]+filter[1500]+filter[1501]+filter[1502]+filter[1503]+filter[1504]+filter[1505]+filter[1506]+filter[1507]+filter[1508]+filter[1509]+filter[1510]+filter[1511]+filter[1512]+filter[1513]+filter[1514]+filter[1515]+filter[1516]+filter[1517]+filter[1518]+filter[1519]+filter[1520]+filter[1521]+filter[1522]+filter[1523]+filter[1524]+filter[1525]+filter[1526]+filter[1527]+filter[1528]+filter[1529]+filter[1530]+filter[1531]+filter[1532]+filter[1533]+filter[1534]+filter[1535]+filter[1536]+filter[1537]+filter[1538]+filter[1539]+filter[1540]+filter[1541]+filter[1542]+filter[1543]+filter[1544]+filter[1545]+filter[1546]+filter[1547]+filter[1548]+filter[1549]+filter[1550]+filter[1551]+filter[1552]+filter[1553]+filter[1554]+filter[1555]+filter[1556]+filter[1557]+filter[1558]+filter[1559]+filter[1560]+filter[1561]+filter[1562]+filter[1563]+filter[1564]+filter[1565]+filter[1566]+filter[1567]+filter[1568]+filter[1569]+filter[1570]+filter[1571]+filter[1572]+filter[1573]+filter[1574]+filter[1575]+filter[1576]+filter[1577]+filter[1578]+filter[1579]+filter[1580]+filter[1581]+filter[1582]+filter[1583]+filter[1584]+filter[1585]+filter[1586]+filter[1587]+filter[1588]+filter[1589]+filter[1590]+filter[1591]+filter[1592]+filter[1593]+filter[1594]+filter[1595]+filter[1596]+filter[1597]+filter[1598]+filter[1599]+filter[1600]+filter[1601]+filter[1602]+filter[1603]+filter[1604]+filter[1605]+filter[1606]+filter[1607]+filter[1608]+filter[1609]+filter[1610]+filter[1611]+filter[1612]+filter[1613]+filter[1614]+filter[1615]+filter[1616]+filter[1617]+filter[1618]+filter[1619]+filter[1620]+filter[1621]+filter[1622]+filter[1623]+filter[1624]+filter[1625]+filter[1626]+filter[1627]+filter[1628]+filter[1629]+filter[1630]+filter[1631]+filter[1632]+filter[1633]+filter[1634]+filter[1635]+filter[1636]+filter[1637]+filter[1638]+filter[1639]+filter[1640]+filter[1641]+filter[1642]+filter[1643]+filter[1644]+filter[1645]+filter[1646]+filter[1647]+filter[1648]+filter[1649]+filter[1650]+filter[1651]+filter[1652]+filter[1653]+filter[1654]+filter[1655]+filter[1656]+filter[1657]+filter[1658]+filter[1659]+filter[1660]+filter[1661]+filter[1662]+filter[1663]+filter[1664]+filter[1665]+filter[1666]+filter[1667]+filter[1668]+filter[1669]+filter[1670]+filter[1671]+filter[1672]+filter[1673]+filter[1674]+filter[1675]+filter[1676]+filter[1677]+filter[1678]+filter[1679]+filter[1680]+filter[1681]+filter[1682]+filter[1683]+filter[1684]+filter[1685]+filter[1686]+filter[1687]+filter[1688]+filter[1689]+filter[1690]+filter[1691]+filter[1692]+filter[1693]+filter[1694]+filter[1695]+filter[1696]+filter[1697]+filter[1698]+filter[1699]+filter[1700]+filter[1701]+filter[1702]+filter[1703]+filter[1704]+filter[1705]+filter[1706]+filter[1707]+filter[1708]+filter[1709]+filter[1710]+filter[1711]+filter[1712]+filter[1713]+filter[1714]+filter[1715]+filter[1716]+filter[1717]+filter[1718]+filter[1719]+filter[1720]+filter[1721]+filter[1722]+filter[1723]+filter[1724]+filter[1725]+filter[1726]+filter[1727]+filter[1728]+filter[1729]+filter[1730]+filter[1731]+filter[1732]+filter[1733]+filter[1734]+filter[1735]+filter[1736]+filter[1737]+filter[1738]+filter[1739]+filter[1740]+filter[1741]+filter[1742]+filter[1743]+filter[1744]+filter[1745]+filter[1746]+filter[1747]+filter[1748]+filter[1749]+filter[1750]+filter[1751]+filter[1752]+filter[1753]+filter[1754]+filter[1755]+filter[1756]+filter[1757]+filter[1758]+filter[1759]+filter[1760]+filter[1761]+filter[1762]+filter[1763]+filter[1764]+filter[1765]+filter[1766]+filter[1767]+filter[1768]+filter[1769]+filter[1770]+filter[1771]+filter[1772]+filter[1773]+filter[1774]+filter[1775]+filter[1776]+filter[1777]+filter[1778]+filter[1779]+filter[1780]+filter[1781]+filter[1782]+filter[1783]+filter[1784]+filter[1785]+filter[1786]+filter[1787]+filter[1788]+filter[1789]+filter[1790]+filter[1791]+filter[1792]+filter[1793]+filter[1794]+filter[1795]+filter[1796]+filter[1797]+filter[1798]+filter[1799]+filter[1800]+filter[1801]+filter[1802]+filter[1803]+filter[1804]+filter[1805]+filter[1806]+filter[1807]+filter[1808]+filter[1809]+filter[1810]+filter[1811]+filter[1812]+filter[1813]+filter[1814]+filter[1815]+filter[1816]+filter[1817]+filter[1818]+filter[1819]+filter[1820]+filter[1821]+filter[1822]+filter[1823]+filter[1824]+filter[1825]+filter[1826]+filter[1827]+filter[1828]+filter[1829]+filter[1830]+filter[1831]+filter[1832]+filter[1833]+filter[1834]+filter[1835]+filter[1836]+filter[1837]+filter[1838]+filter[1839]+filter[1840]+filter[1841]+filter[1842]+filter[1843]+filter[1844]+filter[1845]+filter[1846]+filter[1847]+filter[1848]+filter[1849]+filter[1850]+filter[1851]+filter[1852]+filter[1853]+filter[1854]+filter[1855]+filter[1856]+filter[1857]+filter[1858]+filter[1859]+filter[1860]+filter[1861]+filter[1862]+filter[1863]+filter[1864]+filter[1865]+filter[1866]+filter[1867]+filter[1868]+filter[1869]+filter[1870]+filter[1871]+filter[1872]+filter[1873]+filter[1874]+filter[1875]+filter[1876]+filter[1877]+filter[1878]+filter[1879]+filter[1880]+filter[1881]+filter[1882]+filter[1883]+filter[1884]+filter[1885]+filter[1886]+filter[1887]+filter[1888]+filter[1889]+filter[1890]+filter[1891]+filter[1892]+filter[1893]+filter[1894]+filter[1895]+filter[1896]+filter[1897]+filter[1898]+filter[1899]+filter[1900]+filter[1901]+filter[1902]+filter[1903]+filter[1904]+filter[1905]+filter[1906]+filter[1907]+filter[1908]+filter[1909]+filter[1910]+filter[1911]+filter[1912]+filter[1913]+filter[1914]+filter[1915]+filter[1916]+filter[1917]+filter[1918]+filter[1919]+filter[1920]+filter[1921]+filter[1922]+filter[1923]+filter[1924]+filter[1925]+filter[1926]+filter[1927]+filter[1928]+filter[1929]+filter[1930]+filter[1931]+filter[1932]+filter[1933]+filter[1934]+filter[1935]+filter[1936]+filter[1937]+filter[1938]+filter[1939]+filter[1940]+filter[1941]+filter[1942]+filter[1943]+filter[1944]+filter[1945]+filter[1946]+filter[1947]+filter[1948]+filter[1949]+filter[1950]+filter[1951]+filter[1952]+filter[1953]+filter[1954]+filter[1955]+filter[1956]+filter[1957]+filter[1958]+filter[1959]+filter[1960]+filter[1961]+filter[1962]+filter[1963]+filter[1964]+filter[1965]+filter[1966]+filter[1967]+filter[1968]+filter[1969]+filter[1970]+filter[1971]+filter[1972]+filter[1973]+filter[1974]+filter[1975]+filter[1976]+filter[1977]+filter[1978]+filter[1979]+filter[1980]+filter[1981]+filter[1982]+filter[1983]+filter[1984]+filter[1985]+filter[1986]+filter[1987]+filter[1988]+filter[1989]+filter[1990]+filter[1991]+filter[1992]+filter[1993]+filter[1994]+filter[1995]+filter[1996]+filter[1997]+filter[1998]+filter[1999]+filter[2000]+filter[2001]+filter[2002]+filter[2003]+filter[2004]+filter[2005]+filter[2006]+filter[2007]+filter[2008]+filter[2009]+filter[2010]+filter[2011]+filter[2012]+filter[2013]+filter[2014]+filter[2015]+filter[2016]+filter[2017]+filter[2018]+filter[2019]+filter[2020]+filter[2021]+filter[2022]+filter[2023]+filter[2024]+filter[2025]+filter[2026]+filter[2027]+filter[2028]+filter[2029]+filter[2030]+filter[2031]+filter[2032]+filter[2033]+filter[2034]+filter[2035]+filter[2036]+filter[2037]+filter[2038]+filter[2039]+filter[2040]+filter[2041]+filter[2042]+filter[2043]+filter[2044]+filter[2045]+filter[2046]+filter[2047]+filter[2048]+filter[2049]+filter[2050]+filter[2051]+filter[2052]+filter[2053]+filter[2054]+filter[2055]+filter[2056]+filter[2057]+filter[2058]+filter[2059]+filter[2060]+filter[2061]+filter[2062]+filter[2063]+filter[2064]+filter[2065]+filter[2066]+filter[2067]+filter[2068]+filter[2069]+filter[2070]+filter[2071]+filter[2072]+filter[2073]+filter[2074]+filter[2075]+filter[2076]+filter[2077]+filter[2078]+filter[2079]+filter[2080]+filter[2081]+filter[2082]+filter[2083]+filter[2084]+filter[2085]+filter[2086]+filter[2087]+filter[2088]+filter[2089]+filter[2090]+filter[2091]+filter[2092]+filter[2093]+filter[2094]+filter[2095]+filter[2096]+filter[2097]+filter[2098]+filter[2099]+filter[2100]+filter[2101]+filter[2102]+filter[2103]+filter[2104]+filter[2105]+filter[2106]+filter[2107]+filter[2108]+filter[2109]+filter[2110]+filter[2111]+filter[2112]+filter[2113]+filter[2114]+filter[2115]+filter[2116]+filter[2117]+filter[2118]+filter[2119]+filter[2120]+filter[2121]+filter[2122]+filter[2123]+filter[2124]+filter[2125]+filter[2126]+filter[2127]+filter[2128]+filter[2129]+filter[2130]+filter[2131]+filter[2132]+filter[2133]+filter[2134]+filter[2135]+filter[2136]+filter[2137]+filter[2138]+filter[2139]+filter[2140]+filter[2141]+filter[2142]+filter[2143]+filter[2144]+filter[2145]+filter[2146]+filter[2147]+filter[2148]+filter[2149]+filter[2150]+filter[2151]+filter[2152]+filter[2153]+filter[2154]+filter[2155]+filter[2156]+filter[2157]+filter[2158]+filter[2159]+filter[2160]+filter[2161]+filter[2162]+filter[2163]+filter[2164]+filter[2165]+filter[2166]+filter[2167]+filter[2168]+filter[2169]+filter[2170]+filter[2171]+filter[2172]+filter[2173]+filter[2174]+filter[2175]+filter[2176]+filter[2177]+filter[2178]+filter[2179]+filter[2180]+filter[2181]+filter[2182]+filter[2183]+filter[2184]+filter[2185]+filter[2186]+filter[2187]+filter[2188]+filter[2189]+filter[2190]+filter[2191]+filter[2192]+filter[2193]+filter[2194]+filter[2195]+filter[2196]+filter[2197]+filter[2198]+filter[2199]+filter[2200]+filter[2201]+filter[2202]+filter[2203]+filter[2204]+filter[2205]+filter[2206]+filter[2207]+filter[2208]+filter[2209]+filter[2210]+filter[2211]+filter[2212]+filter[2213]+filter[2214]+filter[2215]+filter[2216]+filter[2217]+filter[2218]+filter[2219]+filter[2220]+filter[2221]+filter[2222]+filter[2223]+filter[2224]+filter[2225]+filter[2226]+filter[2227]+filter[2228]+filter[2229]+filter[2230]+filter[2231]+filter[2232]+filter[2233]+filter[2234]+filter[2235]+filter[2236]+filter[2237]+filter[2238]+filter[2239]+filter[2240]+filter[2241]+filter[2242]+filter[2243]+filter[2244]+filter[2245]+filter[2246]+filter[2247]+filter[2248]+filter[2249]+filter[2250]+filter[2251]+filter[2252]+filter[2253]+filter[2254]+filter[2255]+filter[2256]+filter[2257]+filter[2258]+filter[2259]+filter[2260]+filter[2261]+filter[2262]+filter[2263]+filter[2264]+filter[2265]+filter[2266]+filter[2267]+filter[2268]+filter[2269]+filter[2270]+filter[2271]+filter[2272]+filter[2273]+filter[2274]+filter[2275]+filter[2276]+filter[2277]+filter[2278]+filter[2279]+filter[2280]+filter[2281]+filter[2282]+filter[2283]+filter[2284]+filter[2285]+filter[2286]+filter[2287]+filter[2288]+filter[2289]+filter[2290]+filter[2291]+filter[2292]+filter[2293]+filter[2294]+filter[2295]+filter[2296]+filter[2297]+filter[2298]+filter[2299]+filter[2300]+filter[2301]+filter[2302]+filter[2303]+filter[2304]+filter[2305]+filter[2306]+filter[2307]+filter[2308]+filter[2309]+filter[2310]+filter[2311]+filter[2312]+filter[2313]+filter[2314]+filter[2315]+filter[2316]+filter[2317]+filter[2318]+filter[2319]+filter[2320]+filter[2321]+filter[2322]+filter[2323]+filter[2324]+filter[2325]+filter[2326]+filter[2327]+filter[2328]+filter[2329]+filter[2330]+filter[2331]+filter[2332]+filter[2333]+filter[2334]+filter[2335]+filter[2336]+filter[2337]+filter[2338]+filter[2339]+filter[2340]+filter[2341]+filter[2342]+filter[2343]+filter[2344]+filter[2345]+filter[2346]+filter[2347]+filter[2348]+filter[2349]+filter[2350]+filter[2351]+filter[2352]+filter[2353]+filter[2354]+filter[2355]+filter[2356]+filter[2357]+filter[2358]+filter[2359]+filter[2360]+filter[2361]+filter[2362]+filter[2363]+filter[2364]+filter[2365]+filter[2366]+filter[2367]+filter[2368]+filter[2369]+filter[2370]+filter[2371]+filter[2372]+filter[2373]+filter[2374]+filter[2375]+filter[2376]+filter[2377]+filter[2378]+filter[2379]+filter[2380]+filter[2381]+filter[2382]+filter[2383]+filter[2384]+filter[2385]+filter[2386]+filter[2387]+filter[2388]+filter[2389]+filter[2390]+filter[2391]+filter[2392]+filter[2393]+filter[2394]+filter[2395]+filter[2396]+filter[2397]+filter[2398]+filter[2399]+filter[2400]+filter[2401]+filter[2402]+filter[2403]+filter[2404]+filter[2405]+filter[2406]+filter[2407]+filter[2408]+filter[2409]+filter[2410]+filter[2411]+filter[2412]+filter[2413]+filter[2414]+filter[2415]+filter[2416]+filter[2417]+filter[2418]+filter[2419]+filter[2420]+filter[2421]+filter[2422]+filter[2423]+filter[2424]+filter[2425]+filter[2426]+filter[2427]+filter[2428]+filter[2429]+filter[2430]+filter[2431]+filter[2432]+filter[2433]+filter[2434]+filter[2435]+filter[2436]+filter[2437]+filter[2438]+filter[2439]+filter[2440]+filter[2441]+filter[2442]+filter[2443]+filter[2444]+filter[2445]+filter[2446]+filter[2447]+filter[2448]+filter[2449]+filter[2450]+filter[2451]+filter[2452]+filter[2453]+filter[2454]+filter[2455]+filter[2456]+filter[2457]+filter[2458]+filter[2459]+filter[2460]+filter[2461]+filter[2462]+filter[2463]+filter[2464]+filter[2465]+filter[2466]+filter[2467]+filter[2468]+filter[2469]+filter[2470]+filter[2471]+filter[2472]+filter[2473]+filter[2474]+filter[2475]+filter[2476]+filter[2477]+filter[2478]+filter[2479]+filter[2480]+filter[2481]+filter[2482]+filter[2483]+filter[2484]+filter[2485]+filter[2486]+filter[2487]+filter[2488]+filter[2489]+filter[2490]+filter[2491]+filter[2492]+filter[2493]+filter[2494]+filter[2495]+filter[2496]+filter[2497]+filter[2498]+filter[2499]+filter[2500]+filter[2501]+filter[2502]+filter[2503]+filter[2504]+filter[2505]+filter[2506]+filter[2507]+filter[2508]+filter[2509]+filter[2510]+filter[2511]+filter[2512]+filter[2513]+filter[2514]+filter[2515]+filter[2516]+filter[2517]+filter[2518]+filter[2519]+filter[2520]+filter[2521]+filter[2522]+filter[2523]+filter[2524]+filter[2525]+filter[2526]+filter[2527]+filter[2528]+filter[2529]+filter[2530]+filter[2531]+filter[2532]+filter[2533]+filter[2534]+filter[2535]+filter[2536]+filter[2537]+filter[2538]+filter[2539]+filter[2540]+filter[2541]+filter[2542]+filter[2543]+filter[2544]+filter[2545]+filter[2546]+filter[2547]+filter[2548]+filter[2549]+filter[2550]+filter[2551]+filter[2552]+filter[2553]+filter[2554]+filter[2555]+filter[2556]+filter[2557]+filter[2558]+filter[2559]+filter[2560]+filter[2561]+filter[2562]+filter[2563]+filter[2564]+filter[2565]+filter[2566]+filter[2567]+filter[2568]+filter[2569]+filter[2570]+filter[2571]+filter[2572]+filter[2573]+filter[2574]+filter[2575]+filter[2576]+filter[2577]+filter[2578]+filter[2579]+filter[2580]+filter[2581]+filter[2582]+filter[2583]+filter[2584]+filter[2585]+filter[2586]+filter[2587]+filter[2588]+filter[2589]+filter[2590]+filter[2591]+filter[2592]+filter[2593]+filter[2594]+filter[2595]+filter[2596]+filter[2597]+filter[2598]+filter[2599]+filter[2600]+filter[2601]+filter[2602]+filter[2603]+filter[2604]+filter[2605]+filter[2606]+filter[2607]+filter[2608]+filter[2609]+filter[2610]+filter[2611]+filter[2612]+filter[2613]+filter[2614]+filter[2615]+filter[2616]+filter[2617]+filter[2618]+filter[2619]+filter[2620]+filter[2621]+filter[2622]+filter[2623]+filter[2624]+filter[2625]+filter[2626]+filter[2627]+filter[2628]+filter[2629]+filter[2630]+filter[2631]+filter[2632]+filter[2633]+filter[2634]+filter[2635]+filter[2636]+filter[2637]+filter[2638]+filter[2639]+filter[2640]+filter[2641]+filter[2642]+filter[2643]+filter[2644]+filter[2645]+filter[2646]+filter[2647]+filter[2648]+filter[2649]+filter[2650]+filter[2651]+filter[2652]+filter[2653]+filter[2654]+filter[2655]+filter[2656]+filter[2657]+filter[2658]+filter[2659]+filter[2660]+filter[2661]+filter[2662]+filter[2663]+filter[2664]+filter[2665]+filter[2666]+filter[2667]+filter[2668]+filter[2669]+filter[2670]+filter[2671]+filter[2672]+filter[2673]+filter[2674]+filter[2675]+filter[2676]+filter[2677]+filter[2678]+filter[2679]+filter[2680]+filter[2681]+filter[2682]+filter[2683]+filter[2684]+filter[2685]+filter[2686]+filter[2687]+filter[2688]+filter[2689]+filter[2690]+filter[2691]+filter[2692]+filter[2693]+filter[2694]+filter[2695]+filter[2696]+filter[2697]+filter[2698]+filter[2699]+filter[2700]+filter[2701]+filter[2702]+filter[2703]+filter[2704]+filter[2705]+filter[2706]+filter[2707]+filter[2708]+filter[2709]+filter[2710]+filter[2711]+filter[2712]+filter[2713]+filter[2714]+filter[2715]+filter[2716]+filter[2717]+filter[2718]+filter[2719]+filter[2720]+filter[2721]+filter[2722]+filter[2723]+filter[2724]+filter[2725]+filter[2726]+filter[2727]+filter[2728]+filter[2729]+filter[2730]+filter[2731]+filter[2732]+filter[2733]+filter[2734]+filter[2735]+filter[2736]+filter[2737]+filter[2738]+filter[2739]+filter[2740]+filter[2741]+filter[2742]+filter[2743]+filter[2744]+filter[2745]+filter[2746]+filter[2747]+filter[2748]+filter[2749]+filter[2750]+filter[2751]+filter[2752]+filter[2753]+filter[2754]+filter[2755]+filter[2756]+filter[2757]+filter[2758]+filter[2759]+filter[2760]+filter[2761]+filter[2762]+filter[2763]+filter[2764]+filter[2765]+filter[2766]+filter[2767]+filter[2768]+filter[2769]+filter[2770]+filter[2771]+filter[2772]+filter[2773]+filter[2774]+filter[2775]+filter[2776]+filter[2777]+filter[2778]+filter[2779]+filter[2780]+filter[2781]+filter[2782]+filter[2783]+filter[2784]+filter[2785]+filter[2786]+filter[2787]+filter[2788]+filter[2789]+filter[2790]+filter[2791]+filter[2792]+filter[2793]+filter[2794]+filter[2795]+filter[2796]+filter[2797]+filter[2798]+filter[2799]+filter[2800]+filter[2801]+filter[2802]+filter[2803]+filter[2804]+filter[2805]+filter[2806]+filter[2807]+filter[2808]+filter[2809]+filter[2810]+filter[2811]+filter[2812]+filter[2813]+filter[2814]+filter[2815]+filter[2816]+filter[2817]+filter[2818]+filter[2819]+filter[2820]+filter[2821]+filter[2822]+filter[2823]+filter[2824]+filter[2825]+filter[2826]+filter[2827]+filter[2828]+filter[2829]+filter[2830]+filter[2831]+filter[2832]+filter[2833]+filter[2834]+filter[2835]+filter[2836]+filter[2837]+filter[2838]+filter[2839]+filter[2840]+filter[2841]+filter[2842]+filter[2843]+filter[2844]+filter[2845]+filter[2846]+filter[2847]+filter[2848]+filter[2849]+filter[2850]+filter[2851]+filter[2852]+filter[2853]+filter[2854]+filter[2855]+filter[2856]+filter[2857]+filter[2858]+filter[2859]+filter[2860]+filter[2861]+filter[2862]+filter[2863]+filter[2864]+filter[2865]+filter[2866]+filter[2867]+filter[2868]+filter[2869]+filter[2870]+filter[2871]+filter[2872]+filter[2873]+filter[2874]+filter[2875]+filter[2876]+filter[2877]+filter[2878]+filter[2879]+filter[2880]+filter[2881]+filter[2882]+filter[2883]+filter[2884]+filter[2885]+filter[2886]+filter[2887]+filter[2888]+filter[2889]+filter[2890]+filter[2891]+filter[2892]+filter[2893]+filter[2894]+filter[2895]+filter[2896]+filter[2897]+filter[2898]+filter[2899]+filter[2900]+filter[2901]+filter[2902]+filter[2903]+filter[2904]+filter[2905]+filter[2906]+filter[2907]+filter[2908]+filter[2909]+filter[2910]+filter[2911]+filter[2912]+filter[2913]+filter[2914]+filter[2915]+filter[2916]+filter[2917]+filter[2918]+filter[2919]+filter[2920]+filter[2921]+filter[2922]+filter[2923]+filter[2924]+filter[2925]+filter[2926]+filter[2927]+filter[2928]+filter[2929]+filter[2930]+filter[2931]+filter[2932]+filter[2933]+filter[2934]+filter[2935]+filter[2936]+filter[2937]+filter[2938]+filter[2939]+filter[2940]+filter[2941]+filter[2942]+filter[2943]+filter[2944]+filter[2945]+filter[2946]+filter[2947]+filter[2948]+filter[2949]+filter[2950]+filter[2951]+filter[2952]+filter[2953]+filter[2954]+filter[2955]+filter[2956]+filter[2957]+filter[2958]+filter[2959]+filter[2960]+filter[2961]+filter[2962]+filter[2963]+filter[2964]+filter[2965]+filter[2966]+filter[2967]+filter[2968]+filter[2969]+filter[2970]+filter[2971]+filter[2972]+filter[2973]+filter[2974]+filter[2975]+filter[2976]+filter[2977]+filter[2978]+filter[2979]+filter[2980]+filter[2981]+filter[2982]+filter[2983]+filter[2984]+filter[2985]+filter[2986]+filter[2987]+filter[2988]+filter[2989]+filter[2990]+filter[2991]+filter[2992]+filter[2993]+filter[2994]+filter[2995]+filter[2996]+filter[2997]+filter[2998]+filter[2999]+filter[3000]+filter[3001]+filter[3002]+filter[3003]+filter[3004]+filter[3005]+filter[3006]+filter[3007]+filter[3008]+filter[3009]+filter[3010]+filter[3011]+filter[3012]+filter[3013]+filter[3014]+filter[3015]+filter[3016]+filter[3017]+filter[3018]+filter[3019]+filter[3020]+filter[3021]+filter[3022]+filter[3023]+filter[3024]+filter[3025]+filter[3026]+filter[3027]+filter[3028]+filter[3029]+filter[3030]+filter[3031]+filter[3032]+filter[3033]+filter[3034]+filter[3035]+filter[3036]+filter[3037]+filter[3038]+filter[3039]+filter[3040]+filter[3041]+filter[3042]+filter[3043]+filter[3044]+filter[3045]+filter[3046]+filter[3047]+filter[3048]+filter[3049]+filter[3050]+filter[3051]+filter[3052]+filter[3053]+filter[3054]+filter[3055]+filter[3056]+filter[3057]+filter[3058]+filter[3059]+filter[3060]+filter[3061]+filter[3062]+filter[3063]+filter[3064]+filter[3065]+filter[3066]+filter[3067]+filter[3068]+filter[3069]+filter[3070]+filter[3071]+filter[3072]+filter[3073]+filter[3074]+filter[3075]+filter[3076]+filter[3077]+filter[3078]+filter[3079]+filter[3080]+filter[3081]+filter[3082]+filter[3083]+filter[3084]+filter[3085]+filter[3086]+filter[3087]+filter[3088]+filter[3089]+filter[3090]+filter[3091]+filter[3092]+filter[3093]+filter[3094]+filter[3095]+filter[3096]+filter[3097]+filter[3098]+filter[3099]+filter[3100]+filter[3101]+filter[3102]+filter[3103]+filter[3104]+filter[3105]+filter[3106]+filter[3107]+filter[3108]+filter[3109]+filter[3110]+filter[3111]+filter[3112]+filter[3113]+filter[3114]+filter[3115]+filter[3116]+filter[3117]+filter[3118]+filter[3119]+filter[3120]+filter[3121]+filter[3122]+filter[3123]+filter[3124]+filter[3125]+filter[3126]+filter[3127]+filter[3128]+filter[3129]+filter[3130]+filter[3131]+filter[3132]+filter[3133]+filter[3134]+filter[3135]+filter[3136]+filter[3137]+filter[3138]+filter[3139]+filter[3140]+filter[3141]+filter[3142]+filter[3143]+filter[3144]+filter[3145]+filter[3146]+filter[3147]+filter[3148]+filter[3149]+filter[3150]+filter[3151]+filter[3152]+filter[3153]+filter[3154]+filter[3155]+filter[3156]+filter[3157]+filter[3158]+filter[3159]+filter[3160]+filter[3161]+filter[3162]+filter[3163]+filter[3164]+filter[3165]+filter[3166]+filter[3167]+filter[3168]+filter[3169]+filter[3170]+filter[3171]+filter[3172]+filter[3173]+filter[3174]+filter[3175]+filter[3176]+filter[3177]+filter[3178]+filter[3179]+filter[3180]+filter[3181]+filter[3182]+filter[3183]+filter[3184]+filter[3185]+filter[3186]+filter[3187]+filter[3188]+filter[3189]+filter[3190]+filter[3191]+filter[3192]+filter[3193]+filter[3194]+filter[3195]+filter[3196]+filter[3197]+filter[3198]+filter[3199]+filter[3200]+filter[3201]+filter[3202]+filter[3203]+filter[3204]+filter[3205]+filter[3206]+filter[3207]+filter[3208]+filter[3209]+filter[3210]+filter[3211]+filter[3212]+filter[3213]+filter[3214]+filter[3215]+filter[3216]+filter[3217]+filter[3218]+filter[3219]+filter[3220]+filter[3221]+filter[3222]+filter[3223]+filter[3224]+filter[3225]+filter[3226]+filter[3227]+filter[3228]+filter[3229]+filter[3230]+filter[3231]+filter[3232]+filter[3233]+filter[3234]+filter[3235]+filter[3236]+filter[3237]+filter[3238]+filter[3239]+filter[3240]+filter[3241]+filter[3242]+filter[3243]+filter[3244]+filter[3245]+filter[3246]+filter[3247]+filter[3248]+filter[3249]+filter[3250]+filter[3251]+filter[3252]+filter[3253]+filter[3254]+filter[3255]+filter[3256]+filter[3257]+filter[3258]+filter[3259]+filter[3260]+filter[3261]+filter[3262]+filter[3263]+filter[3264]+filter[3265]+filter[3266]+filter[3267]+filter[3268]+filter[3269]+filter[3270]+filter[3271]+filter[3272]+filter[3273]+filter[3274]+filter[3275]+filter[3276]+filter[3277]+filter[3278]+filter[3279]+filter[3280]+filter[3281]+filter[3282]+filter[3283]+filter[3284]+filter[3285]+filter[3286]+filter[3287]+filter[3288]+filter[3289]+filter[3290]+filter[3291]+filter[3292]+filter[3293]+filter[3294]+filter[3295]+filter[3296]+filter[3297]+filter[3298]+filter[3299]+filter[3300]+filter[3301]+filter[3302]+filter[3303]+filter[3304]+filter[3305]+filter[3306]+filter[3307]+filter[3308]+filter[3309]+filter[3310]+filter[3311]+filter[3312]+filter[3313]+filter[3314]+filter[3315]+filter[3316]+filter[3317]+filter[3318]+filter[3319]+filter[3320]+filter[3321]+filter[3322]+filter[3323]+filter[3324]+filter[3325]+filter[3326]+filter[3327]+filter[3328]+filter[3329]+filter[3330]+filter[3331]+filter[3332]+filter[3333]+filter[3334]+filter[3335]+filter[3336]+filter[3337]+filter[3338]+filter[3339]+filter[3340]+filter[3341]+filter[3342]+filter[3343]+filter[3344]+filter[3345]+filter[3346]+filter[3347]+filter[3348]+filter[3349]+filter[3350]+filter[3351]+filter[3352]+filter[3353]+filter[3354]+filter[3355]+filter[3356]+filter[3357]+filter[3358]+filter[3359]+filter[3360]+filter[3361]+filter[3362]+filter[3363]+filter[3364]+filter[3365]+filter[3366]+filter[3367]+filter[3368]+filter[3369]+filter[3370]+filter[3371]+filter[3372]+filter[3373]+filter[3374]+filter[3375]+filter[3376]+filter[3377]+filter[3378]+filter[3379]+filter[3380]+filter[3381]+filter[3382]+filter[3383]+filter[3384]+filter[3385]+filter[3386]+filter[3387]+filter[3388]+filter[3389]+filter[3390]+filter[3391]+filter[3392]+filter[3393]+filter[3394]+filter[3395]+filter[3396]+filter[3397]+filter[3398]+filter[3399]+filter[3400]+filter[3401]+filter[3402]+filter[3403]+filter[3404]+filter[3405]+filter[3406]+filter[3407]+filter[3408]+filter[3409]+filter[3410]+filter[3411]+filter[3412]+filter[3413]+filter[3414]+filter[3415]+filter[3416]+filter[3417]+filter[3418]+filter[3419]+filter[3420]+filter[3421]+filter[3422]+filter[3423]+filter[3424]+filter[3425]+filter[3426]+filter[3427]+filter[3428]+filter[3429]+filter[3430]+filter[3431]+filter[3432]+filter[3433]+filter[3434]+filter[3435]+filter[3436]+filter[3437]+filter[3438]+filter[3439]+filter[3440]+filter[3441]+filter[3442]+filter[3443]+filter[3444]+filter[3445]+filter[3446]+filter[3447]+filter[3448]+filter[3449]+filter[3450]+filter[3451]+filter[3452]+filter[3453]+filter[3454]+filter[3455]+filter[3456]+filter[3457]+filter[3458]+filter[3459]+filter[3460]+filter[3461]+filter[3462]+filter[3463]+filter[3464]+filter[3465]+filter[3466]+filter[3467]+filter[3468]+filter[3469]+filter[3470]+filter[3471]+filter[3472]+filter[3473]+filter[3474]+filter[3475]+filter[3476]+filter[3477]+filter[3478]+filter[3479]+filter[3480]+filter[3481]+filter[3482]+filter[3483]+filter[3484]+filter[3485]+filter[3486]+filter[3487]+filter[3488]+filter[3489]+filter[3490]+filter[3491]+filter[3492]+filter[3493]+filter[3494]+filter[3495]+filter[3496]+filter[3497]+filter[3498]+filter[3499]+filter[3500]+filter[3501]+filter[3502]+filter[3503]+filter[3504]+filter[3505]+filter[3506]+filter[3507]+filter[3508]+filter[3509]+filter[3510]+filter[3511]+filter[3512]+filter[3513]+filter[3514]+filter[3515]+filter[3516]+filter[3517]+filter[3518]+filter[3519]+filter[3520]+filter[3521]+filter[3522]+filter[3523]+filter[3524]+filter[3525]+filter[3526]+filter[3527]+filter[3528]+filter[3529]+filter[3530]+filter[3531]+filter[3532]+filter[3533]+filter[3534]+filter[3535]+filter[3536]+filter[3537]+filter[3538]+filter[3539]+filter[3540]+filter[3541]+filter[3542]+filter[3543]+filter[3544]+filter[3545]+filter[3546]+filter[3547]+filter[3548]+filter[3549]+filter[3550]+filter[3551]+filter[3552]+filter[3553]+filter[3554]+filter[3555]+filter[3556]+filter[3557]+filter[3558]+filter[3559]+filter[3560]+filter[3561]+filter[3562]+filter[3563]+filter[3564]+filter[3565]+filter[3566]+filter[3567]+filter[3568]+filter[3569]+filter[3570]+filter[3571]+filter[3572]+filter[3573]+filter[3574]+filter[3575]+filter[3576]+filter[3577]+filter[3578]+filter[3579]+filter[3580]+filter[3581]+filter[3582]+filter[3583]+filter[3584]+filter[3585]+filter[3586]+filter[3587]+filter[3588]+filter[3589]+filter[3590]+filter[3591]+filter[3592]+filter[3593]+filter[3594]+filter[3595]+filter[3596]+filter[3597]+filter[3598]+filter[3599]+filter[3600]+filter[3601]+filter[3602]+filter[3603]+filter[3604]+filter[3605]+filter[3606]+filter[3607]+filter[3608]+filter[3609]+filter[3610]+filter[3611]+filter[3612]+filter[3613]+filter[3614]+filter[3615]+filter[3616]+filter[3617]+filter[3618]+filter[3619]+filter[3620]+filter[3621]+filter[3622]+filter[3623]+filter[3624]+filter[3625]+filter[3626]+filter[3627]+filter[3628]+filter[3629]+filter[3630]+filter[3631]+filter[3632]+filter[3633]+filter[3634]+filter[3635]+filter[3636]+filter[3637]+filter[3638]+filter[3639]+filter[3640]+filter[3641]+filter[3642]+filter[3643]+filter[3644]+filter[3645]+filter[3646]+filter[3647]+filter[3648]+filter[3649]+filter[3650]+filter[3651]+filter[3652]+filter[3653]+filter[3654]+filter[3655]+filter[3656]+filter[3657]+filter[3658]+filter[3659]+filter[3660]+filter[3661]+filter[3662]+filter[3663]+filter[3664]+filter[3665]+filter[3666]+filter[3667]+filter[3668]+filter[3669]+filter[3670]+filter[3671]+filter[3672]+filter[3673]+filter[3674]+filter[3675]+filter[3676]+filter[3677]+filter[3678]+filter[3679]+filter[3680]+filter[3681]+filter[3682]+filter[3683]+filter[3684]+filter[3685]+filter[3686]+filter[3687]+filter[3688]+filter[3689]+filter[3690]+filter[3691]+filter[3692]+filter[3693]+filter[3694]+filter[3695]+filter[3696]+filter[3697]+filter[3698]+filter[3699]+filter[3700]+filter[3701]+filter[3702]+filter[3703]+filter[3704]+filter[3705]+filter[3706]+filter[3707]+filter[3708]+filter[3709]+filter[3710]+filter[3711]+filter[3712]+filter[3713]+filter[3714]+filter[3715]+filter[3716]+filter[3717]+filter[3718]+filter[3719]+filter[3720]+filter[3721]+filter[3722]+filter[3723]+filter[3724]+filter[3725]+filter[3726]+filter[3727]+filter[3728]+filter[3729]+filter[3730]+filter[3731]+filter[3732]+filter[3733]+filter[3734]+filter[3735]+filter[3736]+filter[3737]+filter[3738]+filter[3739]+filter[3740]+filter[3741]+filter[3742]+filter[3743]+filter[3744]+filter[3745]+filter[3746]+filter[3747]+filter[3748]+filter[3749]+filter[3750]+filter[3751]+filter[3752]+filter[3753]+filter[3754]+filter[3755]+filter[3756]+filter[3757]+filter[3758]+filter[3759]+filter[3760]+filter[3761]+filter[3762]+filter[3763]+filter[3764]+filter[3765]+filter[3766]+filter[3767]+filter[3768]+filter[3769]+filter[3770]+filter[3771]+filter[3772]+filter[3773]+filter[3774]+filter[3775]+filter[3776]+filter[3777]+filter[3778]+filter[3779]+filter[3780]+filter[3781]+filter[3782]+filter[3783]+filter[3784]+filter[3785]+filter[3786]+filter[3787]+filter[3788]+filter[3789]+filter[3790]+filter[3791]+filter[3792]+filter[3793]+filter[3794]+filter[3795]+filter[3796]+filter[3797]+filter[3798]+filter[3799]+filter[3800]+filter[3801]+filter[3802]+filter[3803]+filter[3804]+filter[3805]+filter[3806]+filter[3807]+filter[3808]+filter[3809]+filter[3810]+filter[3811]+filter[3812]+filter[3813]+filter[3814]+filter[3815]+filter[3816]+filter[3817]+filter[3818]+filter[3819]+filter[3820]+filter[3821]+filter[3822]+filter[3823]+filter[3824]+filter[3825]+filter[3826]+filter[3827]+filter[3828]+filter[3829]+filter[3830]+filter[3831]+filter[3832]+filter[3833]+filter[3834]+filter[3835]+filter[3836]+filter[3837]+filter[3838]+filter[3839]+filter[3840]+filter[3841]+filter[3842]+filter[3843]+filter[3844]+filter[3845]+filter[3846]+filter[3847]+filter[3848]+filter[3849]+filter[3850]+filter[3851]+filter[3852]+filter[3853]+filter[3854]+filter[3855]+filter[3856]+filter[3857]+filter[3858]+filter[3859]+filter[3860]+filter[3861]+filter[3862]+filter[3863]+filter[3864]+filter[3865]+filter[3866]+filter[3867]+filter[3868]+filter[3869]+filter[3870]+filter[3871]+filter[3872]+filter[3873]+filter[3874]+filter[3875]+filter[3876]+filter[3877]+filter[3878]+filter[3879]+filter[3880]+filter[3881]+filter[3882]+filter[3883]+filter[3884]+filter[3885]+filter[3886]+filter[3887]+filter[3888]+filter[3889]+filter[3890]+filter[3891]+filter[3892]+filter[3893]+filter[3894]+filter[3895]+filter[3896]+filter[3897]+filter[3898]+filter[3899]+filter[3900]+filter[3901]+filter[3902]+filter[3903]+filter[3904]+filter[3905]+filter[3906]+filter[3907]+filter[3908]+filter[3909]+filter[3910]+filter[3911]+filter[3912]+filter[3913]+filter[3914]+filter[3915]+filter[3916]+filter[3917]+filter[3918]+filter[3919]+filter[3920]+filter[3921]+filter[3922]+filter[3923]+filter[3924]+filter[3925]+filter[3926]+filter[3927]+filter[3928]+filter[3929]+filter[3930]+filter[3931]+filter[3932]+filter[3933]+filter[3934]+filter[3935]+filter[3936]+filter[3937]+filter[3938]+filter[3939]+filter[3940]+filter[3941]+filter[3942]+filter[3943]+filter[3944]+filter[3945]+filter[3946]+filter[3947]+filter[3948]+filter[3949]+filter[3950]+filter[3951]+filter[3952]+filter[3953]+filter[3954]+filter[3955]+filter[3956]+filter[3957]+filter[3958]+filter[3959]+filter[3960]+filter[3961]+filter[3962]+filter[3963]+filter[3964]+filter[3965]+filter[3966]+filter[3967]+filter[3968]+filter[3969]+filter[3970]+filter[3971]+filter[3972]+filter[3973]+filter[3974]+filter[3975]+filter[3976]+filter[3977]+filter[3978]+filter[3979]+filter[3980]+filter[3981]+filter[3982]+filter[3983]+filter[3984]+filter[3985]+filter[3986]+filter[3987]+filter[3988]+filter[3989]+filter[3990]+filter[3991]+filter[3992]+filter[3993]+filter[3994]+filter[3995]+filter[3996]+filter[3997]+filter[3998]+filter[3999]+filter[4000]+filter[4001]+filter[4002]+filter[4003]+filter[4004]+filter[4005]+filter[4006]+filter[4007]+filter[4008]+filter[4009]+filter[4010]+filter[4011]+filter[4012]+filter[4013]+filter[4014]+filter[4015]+filter[4016]+filter[4017]+filter[4018]+filter[4019]+filter[4020]+filter[4021]+filter[4022]+filter[4023]+filter[4024]+filter[4025]+filter[4026]+filter[4027]+filter[4028]+filter[4029]+filter[4030]+filter[4031]+filter[4032]+filter[4033]+filter[4034]+filter[4035]+filter[4036]+filter[4037]+filter[4038]+filter[4039]+filter[4040]+filter[4041]+filter[4042]+filter[4043]+filter[4044]+filter[4045]+filter[4046]+filter[4047]+filter[4048]+filter[4049]+filter[4050]+filter[4051]+filter[4052]+filter[4053]+filter[4054]+filter[4055]+filter[4056]+filter[4057]+filter[4058]+filter[4059]+filter[4060]+filter[4061]+filter[4062]+filter[4063]+filter[4064]+filter[4065]+filter[4066]+filter[4067]+filter[4068]+filter[4069]+filter[4070]+filter[4071]+filter[4072]+filter[4073]+filter[4074]+filter[4075]+filter[4076]+filter[4077]+filter[4078]+filter[4079]+filter[4080]+filter[4081]+filter[4082]+filter[4083]+filter[4084]+filter[4085]+filter[4086]+filter[4087]+filter[4088]+filter[4089]+filter[4090]+filter[4091]+filter[4092]+filter[4093]+filter[4094]+filter[4095]+filter[4096]+filter[4097]+filter[4098]+filter[4099]+filter[4100]+filter[4101]+filter[4102]+filter[4103]+filter[4104]+filter[4105]+filter[4106]+filter[4107]+filter[4108]+filter[4109]+filter[4110]+filter[4111]+filter[4112]+filter[4113]+filter[4114]+filter[4115]+filter[4116]+filter[4117]+filter[4118]+filter[4119]+filter[4120]+filter[4121]+filter[4122]+filter[4123]+filter[4124]+filter[4125]+filter[4126]+filter[4127]+filter[4128]+filter[4129]+filter[4130]+filter[4131]+filter[4132]+filter[4133]+filter[4134]+filter[4135]+filter[4136]+filter[4137]+filter[4138]+filter[4139]+filter[4140]+filter[4141]+filter[4142]+filter[4143]+filter[4144]+filter[4145]+filter[4146]+filter[4147]+filter[4148]+filter[4149]+filter[4150]+filter[4151]+filter[4152]+filter[4153]+filter[4154]+filter[4155]+filter[4156]+filter[4157]+filter[4158]+filter[4159]+filter[4160]+filter[4161]+filter[4162]+filter[4163]+filter[4164]+filter[4165]+filter[4166]+filter[4167]+filter[4168]+filter[4169]+filter[4170]+filter[4171]+filter[4172]+filter[4173]+filter[4174]+filter[4175]+filter[4176]+filter[4177]+filter[4178]+filter[4179]+filter[4180]+filter[4181]+filter[4182]+filter[4183]+filter[4184]+filter[4185]+filter[4186]+filter[4187]+filter[4188]+filter[4189]+filter[4190]+filter[4191]+filter[4192]+filter[4193]+filter[4194]+filter[4195]+filter[4196]+filter[4197]+filter[4198]+filter[4199]+filter[4200]+filter[4201]+filter[4202]+filter[4203]+filter[4204]+filter[4205]+filter[4206]+filter[4207]+filter[4208]+filter[4209]+filter[4210]+filter[4211]+filter[4212]+filter[4213]+filter[4214]+filter[4215]+filter[4216]+filter[4217]+filter[4218]+filter[4219]+filter[4220]+filter[4221]+filter[4222]+filter[4223]+filter[4224]+filter[4225]+filter[4226]+filter[4227]+filter[4228]+filter[4229]+filter[4230]+filter[4231]+filter[4232]+filter[4233]+filter[4234]+filter[4235]+filter[4236]+filter[4237]+filter[4238]+filter[4239]+filter[4240]+filter[4241]+filter[4242]+filter[4243]+filter[4244]+filter[4245]+filter[4246]+filter[4247]+filter[4248]+filter[4249]+filter[4250]+filter[4251]+filter[4252]+filter[4253]+filter[4254]+filter[4255]+filter[4256]+filter[4257]+filter[4258]+filter[4259]+filter[4260]+filter[4261]+filter[4262]+filter[4263]+filter[4264]+filter[4265]+filter[4266]+filter[4267]+filter[4268]+filter[4269]+filter[4270]+filter[4271]+filter[4272]+filter[4273]+filter[4274]+filter[4275]+filter[4276]+filter[4277]+filter[4278]+filter[4279]+filter[4280]+filter[4281]+filter[4282]+filter[4283]+filter[4284]+filter[4285]+filter[4286]+filter[4287]+filter[4288]+filter[4289]+filter[4290]+filter[4291]+filter[4292]+filter[4293]+filter[4294]+filter[4295]+filter[4296]+filter[4297]+filter[4298]+filter[4299]+filter[4300]+filter[4301]+filter[4302]+filter[4303]+filter[4304]+filter[4305]+filter[4306]+filter[4307]+filter[4308]+filter[4309]+filter[4310]+filter[4311]+filter[4312]+filter[4313]+filter[4314]+filter[4315]+filter[4316]+filter[4317]+filter[4318]+filter[4319]+filter[4320]+filter[4321]+filter[4322]+filter[4323]+filter[4324]+filter[4325]+filter[4326]+filter[4327]+filter[4328]+filter[4329]+filter[4330]+filter[4331]+filter[4332]+filter[4333]+filter[4334]+filter[4335]+filter[4336]+filter[4337]+filter[4338]+filter[4339]+filter[4340]+filter[4341]+filter[4342]+filter[4343]+filter[4344]+filter[4345]+filter[4346]+filter[4347]+filter[4348]+filter[4349]+filter[4350]+filter[4351]+filter[4352]+filter[4353]+filter[4354]+filter[4355]+filter[4356]+filter[4357]+filter[4358]+filter[4359]+filter[4360]+filter[4361]+filter[4362]+filter[4363]+filter[4364]+filter[4365]+filter[4366]+filter[4367]+filter[4368]+filter[4369]+filter[4370]+filter[4371]+filter[4372]+filter[4373]+filter[4374]+filter[4375]+filter[4376]+filter[4377]+filter[4378]+filter[4379]+filter[4380]+filter[4381]+filter[4382]+filter[4383]+filter[4384]+filter[4385]+filter[4386]+filter[4387]+filter[4388]+filter[4389]+filter[4390]+filter[4391]+filter[4392]+filter[4393]+filter[4394]+filter[4395]+filter[4396]+filter[4397]+filter[4398]+filter[4399]+filter[4400]+filter[4401]+filter[4402]+filter[4403]+filter[4404]+filter[4405]+filter[4406]+filter[4407]+filter[4408]+filter[4409]+filter[4410]+filter[4411]+filter[4412]+filter[4413]+filter[4414]+filter[4415]+filter[4416]+filter[4417]+filter[4418]+filter[4419]+filter[4420]+filter[4421]+filter[4422]+filter[4423]+filter[4424]+filter[4425]+filter[4426]+filter[4427]+filter[4428]+filter[4429]+filter[4430]+filter[4431]+filter[4432]+filter[4433]+filter[4434]+filter[4435]+filter[4436]+filter[4437]+filter[4438]+filter[4439]+filter[4440]+filter[4441]+filter[4442]+filter[4443]+filter[4444]+filter[4445]+filter[4446]+filter[4447]+filter[4448]+filter[4449]+filter[4450]+filter[4451]+filter[4452]+filter[4453]+filter[4454]+filter[4455]+filter[4456]+filter[4457]+filter[4458]+filter[4459]+filter[4460]+filter[4461]+filter[4462]+filter[4463]+filter[4464]+filter[4465]+filter[4466]+filter[4467]+filter[4468]+filter[4469]+filter[4470]+filter[4471]+filter[4472]+filter[4473]+filter[4474]+filter[4475]+filter[4476]+filter[4477]+filter[4478]+filter[4479]+filter[4480]+filter[4481]+filter[4482]+filter[4483]+filter[4484]+filter[4485]+filter[4486]+filter[4487]+filter[4488]+filter[4489]+filter[4490]+filter[4491]+filter[4492]+filter[4493]+filter[4494]+filter[4495]+filter[4496]+filter[4497]+filter[4498]+filter[4499]+filter[4500]+filter[4501]+filter[4502]+filter[4503]+filter[4504]+filter[4505]+filter[4506]+filter[4507]+filter[4508]+filter[4509]+filter[4510]+filter[4511]+filter[4512]+filter[4513]+filter[4514]+filter[4515]+filter[4516]+filter[4517]+filter[4518]+filter[4519]+filter[4520]+filter[4521]+filter[4522]+filter[4523]+filter[4524]+filter[4525]+filter[4526]+filter[4527]+filter[4528]+filter[4529]+filter[4530]+filter[4531]+filter[4532]+filter[4533]+filter[4534]+filter[4535]+filter[4536]+filter[4537]+filter[4538]+filter[4539]+filter[4540]+filter[4541]+filter[4542]+filter[4543]+filter[4544]+filter[4545]+filter[4546]+filter[4547]+filter[4548]+filter[4549]+filter[4550]+filter[4551]+filter[4552]+filter[4553]+filter[4554]+filter[4555]+filter[4556]+filter[4557]+filter[4558]+filter[4559]+filter[4560]+filter[4561]+filter[4562]+filter[4563]+filter[4564]+filter[4565]+filter[4566]+filter[4567]+filter[4568]+filter[4569]+filter[4570]+filter[4571]+filter[4572]+filter[4573]+filter[4574]+filter[4575]+filter[4576]+filter[4577]+filter[4578]+filter[4579]+filter[4580]+filter[4581]+filter[4582]+filter[4583]+filter[4584]+filter[4585]+filter[4586]+filter[4587]+filter[4588]+filter[4589]+filter[4590]+filter[4591]+filter[4592]+filter[4593]+filter[4594]+filter[4595]+filter[4596]+filter[4597]+filter[4598]+filter[4599]+filter[4600]+filter[4601]+filter[4602]+filter[4603]+filter[4604]+filter[4605]+filter[4606]+filter[4607]+filter[4608]+filter[4609]+filter[4610]+filter[4611]+filter[4612]+filter[4613]+filter[4614]+filter[4615]+filter[4616]+filter[4617]+filter[4618]+filter[4619]+filter[4620]+filter[4621]+filter[4622]+filter[4623]+filter[4624]+filter[4625]+filter[4626]+filter[4627]+filter[4628]+filter[4629]+filter[4630]+filter[4631]+filter[4632]+filter[4633]+filter[4634]+filter[4635]+filter[4636]+filter[4637]+filter[4638]+filter[4639]+filter[4640]+filter[4641]+filter[4642]+filter[4643]+filter[4644]+filter[4645]+filter[4646]+filter[4647]+filter[4648]+filter[4649]+filter[4650]+filter[4651]+filter[4652]+filter[4653]+filter[4654]+filter[4655]+filter[4656]+filter[4657]+filter[4658]+filter[4659]+filter[4660]+filter[4661]+filter[4662]+filter[4663]+filter[4664]+filter[4665]+filter[4666]+filter[4667]+filter[4668]+filter[4669]+filter[4670]+filter[4671]+filter[4672]+filter[4673]+filter[4674]+filter[4675]+filter[4676]+filter[4677]+filter[4678]+filter[4679]+filter[4680]+filter[4681]+filter[4682]+filter[4683]+filter[4684]+filter[4685]+filter[4686]+filter[4687]+filter[4688]+filter[4689]+filter[4690]+filter[4691]+filter[4692]+filter[4693]+filter[4694]+filter[4695]+filter[4696]+filter[4697]+filter[4698]+filter[4699]+filter[4700]+filter[4701]+filter[4702]+filter[4703]+filter[4704]+filter[4705]+filter[4706]+filter[4707]+filter[4708]+filter[4709]+filter[4710]+filter[4711]+filter[4712]+filter[4713]+filter[4714]+filter[4715]+filter[4716]+filter[4717]+filter[4718]+filter[4719]+filter[4720]+filter[4721]+filter[4722]+filter[4723]+filter[4724]+filter[4725]+filter[4726]+filter[4727]+filter[4728]+filter[4729]+filter[4730]+filter[4731]+filter[4732]+filter[4733]+filter[4734]+filter[4735]+filter[4736]+filter[4737]+filter[4738]+filter[4739]+filter[4740]+filter[4741]+filter[4742]+filter[4743]+filter[4744]+filter[4745]+filter[4746]+filter[4747]+filter[4748]+filter[4749]+filter[4750]+filter[4751]+filter[4752]+filter[4753]+filter[4754]+filter[4755]+filter[4756]+filter[4757]+filter[4758]+filter[4759]+filter[4760]+filter[4761]+filter[4762]+filter[4763]+filter[4764]+filter[4765]+filter[4766]+filter[4767]+filter[4768]+filter[4769]+filter[4770]+filter[4771]+filter[4772]+filter[4773]+filter[4774]+filter[4775]+filter[4776]+filter[4777]+filter[4778]+filter[4779]+filter[4780]+filter[4781]+filter[4782]+filter[4783]+filter[4784]+filter[4785]+filter[4786]+filter[4787]+filter[4788]+filter[4789]+filter[4790]+filter[4791]+filter[4792]+filter[4793]+filter[4794]+filter[4795]+filter[4796]+filter[4797]+filter[4798]+filter[4799]+filter[4800]+filter[4801]+filter[4802]+filter[4803]+filter[4804]+filter[4805]+filter[4806]+filter[4807]+filter[4808]+filter[4809]+filter[4810]+filter[4811]+filter[4812]+filter[4813]+filter[4814]+filter[4815]+filter[4816]+filter[4817]+filter[4818]+filter[4819]+filter[4820]+filter[4821]+filter[4822]+filter[4823]+filter[4824]+filter[4825]+filter[4826]+filter[4827]+filter[4828]+filter[4829]+filter[4830]+filter[4831]+filter[4832]+filter[4833]+filter[4834]+filter[4835]+filter[4836]+filter[4837]+filter[4838]+filter[4839]+filter[4840]+filter[4841]+filter[4842]+filter[4843]+filter[4844]+filter[4845]+filter[4846]+filter[4847]+filter[4848]+filter[4849]+filter[4850]+filter[4851]+filter[4852]+filter[4853]+filter[4854]+filter[4855]+filter[4856]+filter[4857]+filter[4858]+filter[4859]+filter[4860]+filter[4861]+filter[4862]+filter[4863]+filter[4864]+filter[4865]+filter[4866]+filter[4867]+filter[4868]+filter[4869]+filter[4870]+filter[4871]+filter[4872]+filter[4873]+filter[4874]+filter[4875]+filter[4876]+filter[4877]+filter[4878]+filter[4879]+filter[4880]+filter[4881]+filter[4882]+filter[4883]+filter[4884]+filter[4885]+filter[4886]+filter[4887]+filter[4888]+filter[4889]+filter[4890]+filter[4891]+filter[4892]+filter[4893]+filter[4894]+filter[4895]+filter[4896]+filter[4897]+filter[4898]+filter[4899]+filter[4900]+filter[4901]+filter[4902]+filter[4903]+filter[4904]+filter[4905]+filter[4906]+filter[4907]+filter[4908]+filter[4909]+filter[4910]+filter[4911]+filter[4912]+filter[4913]+filter[4914]+filter[4915]+filter[4916]+filter[4917]+filter[4918]+filter[4919]+filter[4920]+filter[4921]+filter[4922]+filter[4923]+filter[4924]+filter[4925]+filter[4926]+filter[4927]+filter[4928]+filter[4929]+filter[4930]+filter[4931]+filter[4932]+filter[4933]+filter[4934]+filter[4935]+filter[4936]+filter[4937]+filter[4938]+filter[4939]+filter[4940]+filter[4941]+filter[4942]+filter[4943]+filter[4944]+filter[4945]+filter[4946]+filter[4947]+filter[4948]+filter[4949]+filter[4950]+filter[4951]+filter[4952]+filter[4953]+filter[4954]+filter[4955]+filter[4956]+filter[4957]+filter[4958]+filter[4959]+filter[4960]+filter[4961]+filter[4962]+filter[4963]+filter[4964]+filter[4965]+filter[4966]+filter[4967]+filter[4968]+filter[4969]+filter[4970]+filter[4971]+filter[4972]+filter[4973]+filter[4974]+filter[4975]+filter[4976]+filter[4977]+filter[4978]+filter[4979]+filter[4980]+filter[4981]+filter[4982]+filter[4983]+filter[4984]+filter[4985]+filter[4986]+filter[4987]+filter[4988]+filter[4989]+filter[4990]+filter[4991]+filter[4992]+filter[4993]+filter[4994]+filter[4995]+filter[4996]+filter[4997]+filter[4998]+filter[4999];
    end
endmodule
